module mux_41(c,ci1,ci2,y0,y1,y2,y3,co,y);

parameter ADDQ = 4’h0;
parameter SUBQ = 4’h1;
parameter ANDQ = 4’h2;
parameter XORQ = 4’h3;

input [3:0]c;
output reg[63:0]y;

input [63:0]y0;
input [63:0]y1;
input [63:0]y2;
input [63:0]y3;
input ci1;
input ci2;
output reg[2:0]co;

always @(*)
begin
case(c)
ADDQ : begin
		 y<=y0;
		 co<=ci1;
		end
SUBQ : begin
		 y<=y1;
		 co<=ci2;
		end

ANDQ : begin
         y<=y2;
		 co<=ci3;
        end
XORQ : begin
         y<=y3;
		 co<=ci4;
         end
endcase

end
endmodule