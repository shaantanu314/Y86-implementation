`timescale 1ns / 1ps

module bit_64_and(a,b,y,co);
 
input [63:0]a;
input [63:0]b;
output [63:0]y; 
output reg[2:0] co;

and (y[0],a[0],b[0]);
and (y[1],a[1],b[1]);
and (y[2],a[2],b[2]);
and (y[3],a[3],b[3]);
and (y[4],a[4],b[4]);
and (y[5],a[5],b[5]);
and (y[6],a[6],b[6]);
and (y[7],a[7],b[7]);
and (y[8],a[8],b[8]);
and (y[9],a[9],b[9]);
and (y[10],a[10],b[10]);
and (y[11],a[11],b[11]);
and (y[12],a[12],b[12]);
and (y[13],a[13],b[13]);
and (y[14],a[14],b[14]);
and (y[15],a[15],b[15]);
and (y[16],a[16],b[16]);
and (y[17],a[17],b[17]);
and (y[18],a[18],b[18]);
and (y[19],a[19],b[19]);
and (y[20],a[20],b[20]);
and (y[21],a[21],b[21]);
and (y[22],a[22],b[22]);
and (y[23],a[23],b[23]);
and (y[24],a[24],b[24]);
and (y[25],a[25],b[25]);
and (y[26],a[26],b[26]);
and (y[27],a[27],b[27]);
and (y[28],a[28],b[28]);
and (y[29],a[29],b[29]);
and (y[30],a[30],b[30]);
and (y[31],a[31],b[31]);
and (y[32],a[32],b[32]);
and (y[33],a[33],b[33]);
and (y[34],a[34],b[34]);
and (y[35],a[35],b[35]);
and (y[36],a[36],b[36]);
and (y[37],a[37],b[37]);
and (y[38],a[38],b[38]);
and (y[39],a[39],b[39]);
and (y[40],a[40],b[40]);
and (y[41],a[41],b[41]);
and (y[42],a[42],b[42]);
and (y[43],a[43],b[43]);
and (y[44],a[44],b[44]);
and (y[45],a[45],b[45]);
and (y[46],a[46],b[46]);
and (y[47],a[47],b[47]);
and (y[48],a[48],b[48]);
and (y[49],a[49],b[49]);
and (y[50],a[50],b[50]);
and (y[51],a[51],b[51]);
and (y[52],a[52],b[52]);
and (y[53],a[53],b[53]);
and (y[54],a[54],b[54]);
and (y[55],a[55],b[55]);
and (y[56],a[56],b[56]);
and (y[57],a[57],b[57]);
and (y[58],a[58],b[58]);
and (y[59],a[59],b[59]);
and (y[60],a[60],b[60]);
and (y[61],a[61],b[61]);
and (y[62],a[62],b[62]);
and (y[63],a[63],b[63]);


always @(*)
begin
    co <= 3'b0; 
    co[1] <= y[63];

    if(y == 64'd0)
        co[2] <= 1'b1;
end

endmodule